module example( input logic a,
                input logic b,
                input logic c,
                output logic y);


assign y = ~a..........

endmodule
